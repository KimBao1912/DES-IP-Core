module Inverse_IP (input logic [63:0] inv_ip_input,
                   output logic [63:0] desc_result);
  assign desc_result = {inv_ip_input[24], inv_ip_input[56], inv_ip_input[16], inv_ip_input[48], inv_ip_input[8], inv_ip_input[40], inv_ip_input[0], inv_ip_input[32], inv_ip_input[25], inv_ip_input[57], inv_ip_input[17], inv_ip_input[49], inv_ip_input[9], inv_ip_input[41], inv_ip_input[1], inv_ip_input[33], inv_ip_input[26], inv_ip_input[58], inv_ip_input[18], inv_ip_input[50], inv_ip_input[10], inv_ip_input[42], inv_ip_input[2], inv_ip_input[34], inv_ip_input[27], inv_ip_input[59], inv_ip_input[19], inv_ip_input[51], inv_ip_input[11], inv_ip_input[43], inv_ip_input[3], inv_ip_input[35], inv_ip_input[28], inv_ip_input[60], inv_ip_input[20], inv_ip_input[52], inv_ip_input[12], inv_ip_input[44], inv_ip_input[4], inv_ip_input[36], inv_ip_input[29], inv_ip_input[61], inv_ip_input[21], inv_ip_input[53], inv_ip_input[13], inv_ip_input[45], inv_ip_input[5], inv_ip_input[37], inv_ip_input[30], inv_ip_input[62], inv_ip_input[22], inv_ip_input[54], inv_ip_input[14], inv_ip_input[46], inv_ip_input[6], inv_ip_input[38], inv_ip_input[31], inv_ip_input[63], inv_ip_input[23], inv_ip_input[55], inv_ip_input[15], inv_ip_input[47], inv_ip_input[7], inv_ip_input[39]};
endmodule
